`include "decode.v"
`include "condlogic.v"

module controller (
	clk,
	reset,
	MulOp,
	Instr,
	MulOp,
	ALUFlags,
	FPUFlags,
	RegSrc,
	RegWrite,
	ImmSrc,
	ALUSrc,
	ALUControl,
	MemWrite,
	MemtoReg,
	PCSrc,
	ResSrc,
	FPUControl
);
	input wire clk;
	input wire reset;
	input wire [7:4] MulOp;
	input wire [31:12] Instr;
	input wire [3:0] ALUFlags;
	input wire [3:0] FPUFlags;
	output wire [1:0] RegSrc;
	output wire RegWrite;
	output wire [1:0] ImmSrc;
	output wire ALUSrc;
	output wire [1:0] ALUControl;
	output wire MemWrite;
	output wire MemtoReg;
	output wire PCSrc;
	output wire ResSrc;
	output wire [1:0] FPUControl;
	wire [1:0] FlagW;
	wire PCS;
	wire RegW;
	wire MemW;
	wire [1:0] FPUFlagW;
	decode dec(
		.Op(Instr[27:26]),
		.Funct(Instr[25:20]),
		.Rd(Instr[15:12]),
		.MulOp(MulOp),
		.FlagW(FlagW),
		.PCS(PCS),
		.RegW(RegW),
		.MemW(MemW),
		.MemtoReg(MemtoReg),
		.ALUSrc(ALUSrc),
		.ImmSrc(ImmSrc),
		.RegSrc(RegSrc),
		.ALUControl(ALUControl),
		.FPUControl(FPUControl),
		.ResSrc(ResSrc),
		.FPUFlagW(FPUFlagW)
	);
	condlogic cl(
		.clk(clk),
		.reset(reset),
		.Cond(Instr[31:28]),
		.ALUFlags(ALUFlags),
		.FPUFlags(FPUFlags),
		.FlagW(FlagW),
		.PCS(PCS),
		.RegW(RegW),
		.MemW(MemW),
		.ResSrc(ResSrc),
		.FPUFlagW(FPUFlagW),
		.PCSrc(PCSrc),
		.RegWrite(RegWrite),
		.MemWrite(MemWrite)
	);
endmodule